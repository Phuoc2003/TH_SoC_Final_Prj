// system_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module system_tb (
	);

	wire        system_inst_clk_bfm_clk_clk;                     // system_inst_clk_bfm:clk -> [system_inst:clk_clk, system_inst_reset_bfm:clk]
	wire  [0:0] system_inst_i2c_0_i2c_serial_bfm_conduit_sda_in; // system_inst_i2c_0_i2c_serial_bfm:sig_sda_in -> system_inst:i2c_0_i2c_serial_sda_in
	wire        system_inst_i2c_0_i2c_serial_sda_oe;             // system_inst:i2c_0_i2c_serial_sda_oe -> system_inst_i2c_0_i2c_serial_bfm:sig_sda_oe
	wire  [0:0] system_inst_i2c_0_i2c_serial_bfm_conduit_scl_in; // system_inst_i2c_0_i2c_serial_bfm:sig_scl_in -> system_inst:i2c_0_i2c_serial_scl_in
	wire        system_inst_i2c_0_i2c_serial_scl_oe;             // system_inst:i2c_0_i2c_serial_scl_oe -> system_inst_i2c_0_i2c_serial_bfm:sig_scl_oe
	wire        system_inst_reset_bfm_reset_reset;               // system_inst_reset_bfm:reset -> system_inst:reset_reset_n

	system system_inst (
		.clk_clk                 (system_inst_clk_bfm_clk_clk),                     //              clk.clk
		.i2c_0_i2c_serial_sda_in (1), // i2c_0_i2c_serial.sda_in
		.i2c_0_i2c_serial_scl_in (1), //                 .scl_in
		.i2c_0_i2c_serial_sda_oe (system_inst_i2c_0_i2c_serial_sda_oe),             //                 .sda_oe
		.i2c_0_i2c_serial_scl_oe (system_inst_i2c_0_i2c_serial_scl_oe),             //                 .scl_oe
		.reset_reset_n           (system_inst_reset_bfm_reset_reset)                //            reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) system_inst_clk_bfm (
		.clk (system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm system_inst_i2c_0_i2c_serial_bfm (
		.sig_scl_in (system_inst_i2c_0_i2c_serial_bfm_conduit_scl_in), // conduit.scl_in
		.sig_scl_oe (system_inst_i2c_0_i2c_serial_scl_oe),             //        .scl_oe
		.sig_sda_in (system_inst_i2c_0_i2c_serial_bfm_conduit_sda_in), //        .sda_in
		.sig_sda_oe (system_inst_i2c_0_i2c_serial_sda_oe)              //        .sda_oe
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) system_inst_reset_bfm (
		.reset (system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
